module shift_reg #(
    parameter DATA_WIDTH = 8
)(
    input wire clk,
    input wire wr_en,
    output reg register[DATA_WIDTH - 1 : 0]
);


endmodule : shift_reg